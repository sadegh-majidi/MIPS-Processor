module control_unit();
